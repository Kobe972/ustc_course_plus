module top(
input		rx,
output	tx);
	assign	tx = rx;
endmodule
